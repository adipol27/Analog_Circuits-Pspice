** Profile: "SCHEMATIC1-anothersim"  [ C:\Users\Or\Desktop\pspicecircuits\0602proj-pspicefiles\schematic1\anothersim.sim ] 

** Creating circuit file "anothersim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../0602proj-pspicefiles/0602proj.lib" 
* From [PSPICE NETLIST] section of C:\Users\Or\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.AC DEC 1000 100Hz 100MegHz
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
